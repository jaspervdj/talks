<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->
<svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:cc="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" xmlns:svg="http://www.w3.org/2000/svg" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape" width="256" height="256" id="svg2" sodipodi:version="0.32" inkscape:version="0.47 r22583" sodipodi:docname="blogger.svg" version="1.0" inkscape:output_extension="org.inkscape.output.svg.inkscape">
  <defs id="defs4">
    <linearGradient inkscape:collect="always" id="linearGradient2555">
      <stop style="stop-color: rgb(255, 255, 255); stop-opacity: 1;" offset="0" id="stop2557"/>
      <stop style="stop-color: rgb(255, 255, 255); stop-opacity: 0;" offset="1" id="stop2559"/>
    </linearGradient>
    <linearGradient inkscape:collect="always" xlink:href="#linearGradient2555" id="linearGradient2449" gradientUnits="userSpaceOnUse" gradientTransform="matrix(-0.5914583,0,0,0.5914584,210.0216,142.2324)" x1="-344.15295" y1="274.711" x2="-395.84943" y2="425.39993"/>
  </defs>
  <sodipodi:namedview id="base" pagecolor="#ffffff" bordercolor="#666666" borderopacity="1.0" inkscape:pageopacity="0.0" inkscape:pageshadow="2" inkscape:zoom="0.24748737" inkscape:cx="150.19857" inkscape:cy="122.62969" inkscape:document-units="px" inkscape:current-layer="layer1" inkscape:window-width="782" inkscape:window-height="674" inkscape:window-x="1" inkscape:window-y="281" showgrid="false" inkscape:window-maximized="0"/>
  <metadata id="metadata7">
    <rdf:RDF>
      <cc:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
        <dc:creator>
          <cc:Agent>
            <dc:title/>
          </cc:Agent>
        </dc:creator>
        <dc:subject>
          <rdf:Bag/>
        </dc:subject>
        <cc:license rdf:resource="http://creativecommons.org/licenses/publicdomain/"/>
        <dc:description/>
        <dc:contributor>
          <cc:Agent>
            <dc:title/>
          </cc:Agent>
        </dc:contributor>
      </cc:Work>
      <cc:License rdf:about="http://creativecommons.org/licenses/publicdomain/">
        <cc:permits rdf:resource="http://creativecommons.org/ns#Reproduction"/>
        <cc:permits rdf:resource="http://creativecommons.org/ns#Distribution"/>
        <cc:permits rdf:resource="http://creativecommons.org/ns#DerivativeWorks"/>
      </cc:License>
    </rdf:RDF>
  </metadata>
  <g inkscape:label="Layer 1" inkscape:groupmode="layer" id="layer1" transform="translate(-373.642,-318.344)">
    <rect inkscape:export-ydpi="7.7063322" inkscape:export-xdpi="7.7063322" inkscape:export-filename="C:\Documents and Settings\Molumen\Desktop\path3511111.png" transform="scale(-1,1)" ry="35.487503" rx="35.487503" y="328.84921" x="-619.14587" height="234.98955" width="235.00784" id="rect1942" style="fill:#f57d00;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:0.87500000000000000;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:0.87500000000000000, 1.75000000000000000;stroke-dashoffset:0;stroke-opacity:1"/>
    <path inkscape:export-ydpi="7.7063322" inkscape:export-xdpi="7.7063322" inkscape:export-filename="C:\Documents and Settings\Molumen\Desktop\path3511111.png" sodipodi:nodetypes="ccccsssc" id="path1950" d="M 557.05665,338.89518 L 446.22721,338.89518 C 416.89033,338.89518 393.27256,362.70492 393.27256,392.28025 L 393.27256,500.40761 C 394.22216,523.49366 397.87485,508.89915 404.82758,483.3329 C 412.90814,453.61975 439.22406,427.65003 471.27219,408.1872 C 495.73352,393.33195 523.11328,383.84595 572.95174,382.94353 C 601.21656,382.43177 598.72124,346.26062 557.05665,338.89518 z" style="opacity:1;fill:url(#linearGradient2449);fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:0.87500000000000000;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:0.87500000000000000, 1.75000000000000000;stroke-dashoffset:0;stroke-opacity:1"/>
    <path style="fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#ffffff;stroke-width:30;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="M 474.28848,392.93948 L 508.3909,392.41491 C 524.00714,392.84658 532.6861,403.91597 532.52493,416.5451 C 534.0387,431.46829 529.83653,448.36648 506.29229,448.01925 L 472.71452,448.01925 C 457.9097,448.16241 446.08833,439.46231 447.00654,422.31536 C 446.27306,408.10943 450.9639,392.73464 474.28848,392.93948 z" id="path3778" sodipodi:nodetypes="ccccccc"/>
    <path style="fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#ffffff;stroke-width:30;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="M 529.37701,508.34471 L 476.91174,508.34471 C 455.04991,508.6252 444.51929,498.65845 445.95723,475.82142 C 446.06053,455.29282 457.96814,449.4313 475.86244,449.06839 L 527.80304,449.06839 C 563.12025,448.12561 559.26294,447.78377 559.80686,476.34598 C 559.58484,497.11094 548.1648,508.18579 529.37701,508.34471 z" id="path3780" sodipodi:nodetypes="ccccccc"/>
    <path style="fill:none;fill-rule:evenodd;stroke:#ffffff;stroke-width:30;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="M 445.95724,480.01797 L 447.00654,417.06966" id="path3782" sodipodi:nodetypes="cc"/>
    <path style="fill:none;fill-rule:evenodd;stroke:#f57d00;stroke-width:25;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="M 476.78254,419.90545 L 506.07336,420.3705" id="path3786" sodipodi:nodetypes="cc"/>
    <path style="fill:none;fill-rule:evenodd;stroke:#f57d00;stroke-width:25;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="M 473.45507,477.18678 L 532.03671,477.18678" id="path3788" sodipodi:nodetypes="cc"/>
  </g>
</svg>